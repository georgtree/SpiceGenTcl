

.dc v1 {time1} 5 0.1
.dc v1 0 5 0.1
.ac dec 10 {f1} 1e6
.ac lin 1000 1 1e6
.sp dec 10 {f1} 1e6
.sp lin 1000 1 1e6
.sp lin 1000 1 1e6 1
.sens v(1, out) ac dec 10 {f1} 1e6
.sens v(1,out ) ac dec 10 1 1e6
.sens v(  1, out) ac dec 10 1 1e6
.sens i(1,out)
.tran 1e-6 1e-3 0.1e-6 uic
.tran 1e-6 {tend} uic
.op
