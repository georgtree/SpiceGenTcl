
.subckt resarr in out PARAMS: rs=2 rt=3
r1 in a r={rs}
r2 a out r={rt}
.ends
.subckt resarr1 in out rs=2 rt=3
r1 in a r={rs}
r2 a out r={rt}
.ends
