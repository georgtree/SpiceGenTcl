

.param u0t={rf+1} vth0=10
.param k1=1e-4 vth0=10 u0t={rf+1 }
.param abv=1 tre= 1k pre=1MEG
