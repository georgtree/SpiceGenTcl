
.subckt resarr in out PARAMS: rs=2 rt=3
r1 in a r={rs}
r2 a out r={rt}
.subckt resarr1 in out rs=2 rt=3
r1 in a r={rs}
r2 a out r={rt}
.subckt resarr2 in out rs=2 rt=3
r1 in a r={rs}
r2 a out r={rt}
.ends
x1 a b resarr2
.ends
x1 a b resarr1
.ends
