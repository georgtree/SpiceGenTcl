

.model resmod r(tc1=1 tc2=2)
.model capmod c tc1=1 tc2=2
.model indmod l( tc1=1 tc2=2)
.model swmod sw(vt=1 vh=0.5 ron=1 roff=1e6 )
.model cswmod csw ( it=1 ih=0.5 ron=1 roff=1e6)
.model diodemod d(is=1e-14 n=1.2 rs=0.01 cjo=1e-9)
.model bjtmod npn (level=1 is=1e-15 bf=200 vaf=100 cje=1e-10)
.model bjtmod1 npn (level=4 is=1e-15 bf=200 vaf=100 cje=1e-10)
.model jfetmod1 njf  level=1 vto=2 beta=1e-3 lambda=1e-4 cgd=1e-12
.model jfetmod2 njf(vto=2 beta=1e-3 lambda=1e-4 cgd=1e-12)
.model jfetmod3 njf(level=2.0 vto=-2 beta=10e-4 rs=1e-4 vbi=1.2)
.model mesfetmod1 nmf(level=1 vto=2 beta=1e-3 lambda=1e-4 cgd=1e-12)
.model mesfetmod2 pmf(vto=-2 beta=1e-3 lambda=1e-4 cgd=1e-12)
.model res3mod r3(tc1=1 tc2=2)
